entity asd is
constant asd : integer := 0;
type asdf is range 0 to 5;
end entity;
