entity asd is
generic (
  type asd;
  constant asd : integer := 0;
);
port ( signal asd : in std_logic(asd) := '0');
constant asd : integer := 0;type asdf is range 0 to 5;
end entity;
