entity asd is
generic (
  type asd;
  constant asd : integer := 0;
);
port ( signal asd : in std_logic(asd) := '0');
constant asd : integer := 0;type asdf is range 0 to 5;
end entity;

architecture asd of gg is
  component asd
    generic( asd : tst := 123);
    port (signal asd:bbb; asd : out fff);
    end component;
impure function test(asd : interger := 1) return integer is
  variable temp : integer := 0;
begin
  return temp;
  end function;
  begin

  end architecture beh;