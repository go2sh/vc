entity asd is
constant �asd : integer := 0;
end entity;
